module		sample1(s, a, b);
	input	a, b;
	output	s;
	assign	s = a & b;
endmodule